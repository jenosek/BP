** Profile: "SCHEMATIC1-frec"  [ C:\Skola\VUT\CubeSat\BP\simulations\PSpice\lp_ant\lp_ant-pspicefiles\schematic1\frec.sim ] 

** Creating circuit file "frec.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\honza\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 1400 1megHz 1GHz
.STEP LIN PARAM c 7pF 14pF 0.1pF 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
